library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package MEMORY_PACK is--Package creation


--The below all statements creates necwssary data vectors which can be used in top module
type RAM_LOC is array(natural range <>) of std_logic_vector;

end package MEMORY_PACK;