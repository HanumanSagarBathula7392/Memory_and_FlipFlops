library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


package MEMORY_PACK is

type RAM_LOC is array(natural range<>) of std_logic_vector;

end package MEMORY_PACK;
